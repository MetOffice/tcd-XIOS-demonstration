netcdf domain_input {
dimensions:
        x = 5 ;
        y = 5 ;
        alt = 1 ;
variables:
        float x(x) ;
                x:standard_name = "projection_x_coordinate" ;
                x:units = "m";
        float y(y) ;
                y:standard_name = "projection_y_coordinate" ;
                y:units = "m";
        float alt(alt) ;
                alt:standard_name = "altitude" ;
                alt:units = "metres";                
        double original_data(alt, y, x) ;
                original_data:long_name = "data values" ;
                original_data:units = "1";

// global attributes:
                :title = "Input data for XIOS output." ;

data:

 x = 303000, 305000, 307000, 309000, 311000 ;

 y = 107000, 109000, 111000, 113000, 115000 ;

 alt = 50 ;

 original_data =  0,  2,  4,  6,  8,
                  2,  4,  6,  8, 10,
                  4,  6,  8, 10, 12,
                  6,  8, 10, 12, 14,
                  8, 10, 12, 14, 16 ;

}
