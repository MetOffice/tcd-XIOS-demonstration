netcdf data_output {
dimensions:
	axis_nbounds = 2 ;
	Two = 2 ;
	ncubedsphere_node = 8 ;
	ncubedsphere_edge = 12 ;
	ncubedsphere_face = 6 ;
	ncubedsphere_vertex = 4 ;
	nmain__domain_undef_id_8_node = 8 ;
	nmain__domain_undef_id_8_edge = 12 ;
	nmain__domain_undef_id_6_node = 8 ;
	time_counter = UNLIMITED ; // (2 currently)
variables:
	int cubedsphere ;
		cubedsphere:cf_role = "mesh_topology" ;
		cubedsphere:long_name = "Topology data of 2D unstructured mesh" ;
		cubedsphere:topology_dimension = 2 ;
		cubedsphere:node_coordinates = "cubedsphere_node_x cubedsphere_node_y" ;
		cubedsphere:edge_coordinates = "cubedsphere_edge_x cubedsphere_edge_y" ;
		cubedsphere:edge_node_connectivity = "cubedsphere_edge_nodes" ;
		cubedsphere:face_edge_connectivity = "cubedsphere_face_edges" ;
		cubedsphere:edge_face_connectivity = "cubedsphere_edge_face_links" ;
		cubedsphere:face_face_connectivity = "cubedsphere_face_links" ;
		cubedsphere:face_coordinates = "cubedsphere_face_x cubedsphere_face_y" ;
		cubedsphere:face_node_connectivity = "cubedsphere_face_nodes" ;
	float cubedsphere_node_x(ncubedsphere_node) ;
		cubedsphere_node_x:standard_name = "longitude" ;
		cubedsphere_node_x:long_name = "Longitude of mesh nodes." ;
		cubedsphere_node_x:units = "degrees_east" ;
	float cubedsphere_node_y(ncubedsphere_node) ;
		cubedsphere_node_y:standard_name = "latitude" ;
		cubedsphere_node_y:long_name = "Latitude of mesh nodes." ;
		cubedsphere_node_y:units = "degrees_north" ;
	float cubedsphere_edge_x(ncubedsphere_edge) ;
		cubedsphere_edge_x:standard_name = "longitude" ;
		cubedsphere_edge_x:long_name = "Characteristic longitude of mesh edges." ;
		cubedsphere_edge_x:units = "degrees_east" ;
	float cubedsphere_edge_y(ncubedsphere_edge) ;
		cubedsphere_edge_y:standard_name = "latitude" ;
		cubedsphere_edge_y:long_name = "Characteristic latitude of mesh edges." ;
		cubedsphere_edge_y:units = "degrees_north" ;
	int cubedsphere_edge_nodes(ncubedsphere_edge, Two) ;
		cubedsphere_edge_nodes:cf_role = "edge_node_connectivity" ;
		cubedsphere_edge_nodes:long_name = "Maps every edge/link to two nodes that it connects." ;
		cubedsphere_edge_nodes:start_index = 0 ;
	float cubedsphere_face_x(ncubedsphere_face) ;
		cubedsphere_face_x:standard_name = "longitude" ;
		cubedsphere_face_x:long_name = "Characteristic longitude of mesh faces." ;
		cubedsphere_face_x:units = "degrees_east" ;
	float cubedsphere_face_y(ncubedsphere_face) ;
		cubedsphere_face_y:standard_name = "latitude" ;
		cubedsphere_face_y:long_name = "Characteristic latitude of mesh faces." ;
		cubedsphere_face_y:units = "degrees_north" ;
	int cubedsphere_face_nodes(ncubedsphere_face, ncubedsphere_vertex) ;
		cubedsphere_face_nodes:cf_role = "face_node_connectivity" ;
		cubedsphere_face_nodes:long_name = "Maps every face to its corner nodes." ;
		cubedsphere_face_nodes:start_index = 0 ;
	int cubedsphere_face_edges(ncubedsphere_face, ncubedsphere_vertex) ;
		cubedsphere_face_edges:cf_role = "face_edge_connectivity" ;
		cubedsphere_face_edges:long_name = "Maps every face to its edges." ;
		cubedsphere_face_edges:start_index = 0 ;
		cubedsphere_face_edges:_FillValue = 999999 ;
	int cubedsphere_edge_face_links(ncubedsphere_edge, Two) ;
		cubedsphere_edge_face_links:cf_role = "edge_face_connectivity" ;
		cubedsphere_edge_face_links:long_name = "neighbor faces for edges" ;
		cubedsphere_edge_face_links:start_index = 0 ;
		cubedsphere_edge_face_links:_FillValue = -999 ;
		cubedsphere_edge_face_links:comment = "missing neighbor faces are indicated using _FillValue" ;
	int cubedsphere_face_links(ncubedsphere_face, ncubedsphere_vertex) ;
		cubedsphere_face_links:cf_role = "face_face_connectivity" ;
		cubedsphere_face_links:long_name = "Indicates which other faces neighbor each face" ;
		cubedsphere_face_links:start_index = 0 ;
		cubedsphere_face_links:_FillValue = 999999 ;
		cubedsphere_face_links:flag_values = -1 ;
		cubedsphere_face_links:flag_meanings = "out_of_mesh" ;
	int main__domain_undef_id_8 ;
		main__domain_undef_id_8:cf_role = "mesh_topology" ;
		main__domain_undef_id_8:long_name = "Topology data of 2D unstructured mesh" ;
		main__domain_undef_id_8:topology_dimension = 2 ;
		main__domain_undef_id_8:node_coordinates = "main__domain_undef_id_8_node_x main__domain_undef_id_8_node_y" ;
		main__domain_undef_id_8:edge_node_connectivity = "main__domain_undef_id_8_edge_nodes" ;
		main__domain_undef_id_8:edge_coordinates = "main__domain_undef_id_8_edge_x main__domain_undef_id_8_edge_y" ;
	float main__domain_undef_id_8_node_x(nmain__domain_undef_id_8_node) ;
		main__domain_undef_id_8_node_x:standard_name = "longitude" ;
		main__domain_undef_id_8_node_x:long_name = "Longitude of mesh nodes." ;
		main__domain_undef_id_8_node_x:units = "degrees_east" ;
	float main__domain_undef_id_8_node_y(nmain__domain_undef_id_8_node) ;
		main__domain_undef_id_8_node_y:standard_name = "latitude" ;
		main__domain_undef_id_8_node_y:long_name = "Latitude of mesh nodes." ;
		main__domain_undef_id_8_node_y:units = "degrees_north" ;
	float main__domain_undef_id_8_edge_x(nmain__domain_undef_id_8_edge) ;
		main__domain_undef_id_8_edge_x:standard_name = "longitude" ;
		main__domain_undef_id_8_edge_x:long_name = "Characteristic longitude of mesh edges." ;
		main__domain_undef_id_8_edge_x:units = "degrees_east" ;
	float main__domain_undef_id_8_edge_y(nmain__domain_undef_id_8_edge) ;
		main__domain_undef_id_8_edge_y:standard_name = "latitude" ;
		main__domain_undef_id_8_edge_y:long_name = "Characteristic latitude of mesh edges." ;
		main__domain_undef_id_8_edge_y:units = "degrees_north" ;
	int main__domain_undef_id_8_edge_nodes(nmain__domain_undef_id_8_edge, Two) ;
		main__domain_undef_id_8_edge_nodes:cf_role = "edge_node_connectivity" ;
		main__domain_undef_id_8_edge_nodes:long_name = "Maps every edge/link to two nodes that it connects." ;
		main__domain_undef_id_8_edge_nodes:start_index = 0 ;
	int main__domain_undef_id_6 ;
		main__domain_undef_id_6:cf_role = "mesh_topology" ;
		main__domain_undef_id_6:long_name = "Topology data of 2D unstructured mesh" ;
		main__domain_undef_id_6:topology_dimension = 2 ;
		main__domain_undef_id_6:node_coordinates = "main__domain_undef_id_6_node_x main__domain_undef_id_6_node_y" ;
	float main__domain_undef_id_6_node_x(nmain__domain_undef_id_6_node) ;
		main__domain_undef_id_6_node_x:standard_name = "longitude" ;
		main__domain_undef_id_6_node_x:long_name = "Longitude of mesh nodes." ;
		main__domain_undef_id_6_node_x:units = "degrees_east" ;
	float main__domain_undef_id_6_node_y(nmain__domain_undef_id_6_node) ;
		main__domain_undef_id_6_node_y:standard_name = "latitude" ;
		main__domain_undef_id_6_node_y:long_name = "Latitude of mesh nodes." ;
		main__domain_undef_id_6_node_y:units = "degrees_north" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-02-02 12:00:00" ;
		time_instant:time_origin = "2022-02-02 12:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-02-02 12:00:00" ;
		time_counter:time_origin = "2022-02-02 12:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	double arbitrary_face_data(time_counter, ncubedsphere_face) ;
		arbitrary_face_data:long_name = "Arbitrary data values" ;
		arbitrary_face_data:units = "1" ;
		arbitrary_face_data:mesh = "cubedsphere" ;
		arbitrary_face_data:location = "face" ;
		arbitrary_face_data:online_operation = "instant" ;
		arbitrary_face_data:interval_operation = "1 h" ;
		arbitrary_face_data:interval_write = "1 h" ;
		arbitrary_face_data:cell_methods = "time: point" ;
		arbitrary_face_data:coordinates = "time_instant cubedsphere_face_y cubedsphere_face_x" ;
	double arbitrary_edge_data(time_counter, nmain__domain_undef_id_8_edge) ;
		arbitrary_edge_data:long_name = "Arbitrary data values" ;
		arbitrary_edge_data:units = "1" ;
		arbitrary_edge_data:mesh = "main__domain_undef_id_8" ;
		arbitrary_edge_data:location = "edge" ;
		arbitrary_edge_data:online_operation = "instant" ;
		arbitrary_edge_data:interval_operation = "1 h" ;
		arbitrary_edge_data:interval_write = "1 h" ;
		arbitrary_edge_data:cell_methods = "time: point" ;
		arbitrary_edge_data:coordinates = "time_instant main__domain_undef_id_8_edge_y main__domain_undef_id_8_edge_x" ;
	double arbitrary_node_data(time_counter, nmain__domain_undef_id_6_node) ;
		arbitrary_node_data:long_name = "Arbitrary data values" ;
		arbitrary_node_data:units = "1" ;
		arbitrary_node_data:mesh = "main__domain_undef_id_6" ;
		arbitrary_node_data:location = "node" ;
		arbitrary_node_data:online_operation = "instant" ;
		arbitrary_node_data:interval_operation = "1 h" ;
		arbitrary_node_data:interval_write = "1 h" ;
		arbitrary_node_data:cell_methods = "time: point" ;
		arbitrary_node_data:coordinates = "time_instant main__domain_undef_id_6_node_y main__domain_undef_id_6_node_x" ;

// global attributes:
		:name = "data_output" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "UGRID" ;
		:timeStamp = "2025-May-07 14:23:04 GMT" ;
		:uuid = "02f24392-2446-494f-a1a7-d482900beb2b" ;
data:

 cubedsphere = _ ;

 cubedsphere_node_x = -45, 45, 135, -135, 45, -45, 135, -135 ;

 cubedsphere_node_y = 35.26439, 35.26439, 35.26439, 35.26439, -35.26439, 
    -35.26439, -35.26439, -35.26439 ;

 cubedsphere_edge_x = 0, -45, 0, 90, 45, 90, 0, 135, 0, -90, -135, -90 ;

 cubedsphere_edge_y = 35.26439, 0, -35.26439, 35.26439, 0, -35.26439, 
    35.26439, 0, -35.26439, 35.26439, 0, -35.26439 ;

 cubedsphere_edge_nodes =
  0, 1,
  5, 0,
  4, 5,
  1, 2,
  4, 1,
  6, 4,
  2, 3,
  6, 2,
  7, 6,
  3, 0,
  7, 3,
  5, 7 ;

 cubedsphere_face_x = 2.754441e-15, 90, -180, -90, 0, 0 ;

 cubedsphere_face_y = -5.508882e-15, -5.508882e-15, -5.508882e-15, 
    -5.508882e-15, 90, -90 ;

 cubedsphere_face_nodes =
  5, 4, 1, 0,
  4, 6, 2, 1,
  7, 3, 2, 6,
  5, 0, 3, 7,
  0, 1, 2, 3,
  5, 7, 6, 4 ;

 cubedsphere_face_edges =
  2, 4, 0, 1,
  5, 7, 3, 4,
  10, 6, 7, 8,
  1, 9, 10, 11,
  0, 3, 6, 9,
  11, 8, 5, 2 ;

 cubedsphere_edge_face_links =
  0, 4,
  0, 3,
  0, 5,
  1, 4,
  0, 1,
  1, 5,
  2, 4,
  1, 2,
  2, 5,
  3, 4,
  2, 3,
  3, 5 ;

 cubedsphere_face_links =
  5, 1, 4, 3,
  5, 2, 4, 0,
  3, 4, 1, 5,
  0, 4, 2, 5,
  0, 1, 2, 3,
  3, 2, 1, 0 ;

 main__domain_undef_id_8 = _ ;

 main__domain_undef_id_8_node_x = -45, 45, 135, -135, 45, -45, 135, -135 ;

 main__domain_undef_id_8_node_y = 35.26439, 35.26439, 35.26439, 35.26439, 
    -35.26439, -35.26439, -35.26439, -35.26439 ;

 main__domain_undef_id_8_edge_x = 0, -45, 0, 90, 45, 90, 0, 135, 0, -90, 
    -135, -90 ;

 main__domain_undef_id_8_edge_y = 35.26439, 0, -35.26439, 35.26439, 0, 
    -35.26439, 35.26439, 0, -35.26439, 35.26439, 0, -35.26439 ;

 main__domain_undef_id_8_edge_nodes =
  0, 1,
  5, 0,
  4, 5,
  1, 2,
  4, 1,
  6, 4,
  2, 3,
  6, 2,
  7, 6,
  3, 0,
  7, 3,
  5, 7 ;

 main__domain_undef_id_6 = _ ;

 main__domain_undef_id_6_node_x = -45, 45, 135, -135, 45, -45, 135, -135 ;

 main__domain_undef_id_6_node_y = 35.26439, 35.26439, 35.26439, 35.26439, 
    -35.26439, -35.26439, -35.26439, -35.26439 ;

 time_instant = 27133200, 27136800 ;

 time_instant_bounds =
  27133200, 27133200,
  27136800, 27136800 ;

 time_counter = 27133200, 27136800 ;

 time_counter_bounds =
  27133200, 27133200,
  27136800, 27136800 ;

 arbitrary_face_data =
  10, 10, 10, 10, 10, 10,
  20, 20, 20, 20, 20, 20 ;

 arbitrary_edge_data =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200 ;

 arbitrary_node_data =
  1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2 ;
}
