netcdf data_output {
dimensions:
	axis_nbounds = 2 ;
	x = 5 ;
	y = 5 ;
	alt = 1 ;
	time_counter = UNLIMITED ; // (1 currently)
variables:
	float x(x) ;
		x:name = "x" ;
		x:standard_name = "projection_x_coordinate" ;
		x:long_name = "x coordinate of projection" ;
		x:units = "m" ;
	float y(y) ;
		y:name = "y" ;
		y:standard_name = "projection_y_coordinate" ;
		y:long_name = "y coordinate of projection" ;
		y:units = "m" ;
	float alt(alt) ;
		alt:name = "alt" ;
		alt:standard_name = "altitude" ;
		alt:units = "metres" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-02-02 12:00:00" ;
		time_instant:time_origin = "2022-02-02 12:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-02-02 12:00:00" ;
		time_counter:time_origin = "2022-02-02 12:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	double forecast_reference_time ;
	        forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "gregorian" ;
		forecast_reference_time:units = "seconds since 2022-02-02 12:00:00" ;
		forecast_reference_time:time_origin = "2022-02-02 12:00:00" ;	
	double original_data(time_counter, alt, y, x) ;
		original_data:long_name = "Arbitrary data values" ;
		original_data:units = "1" ;
		original_data:online_operation = "instant" ;
		original_data:interval_operation = "1 h" ;
		original_data:interval_write = "1 h" ;
		original_data:cell_methods = "time: point" ;
		original_data:coordinates = "time_instant forecast_reference_time" ;

// global attributes:
		:description = "LFRic file format v0.2.0" ;
		:Conventions = "CF-1.6, UGRID" ;
		:timeStamp = "2025-Apr-16 16:24:09 GMT" ;
		:uuid = "faa3e3a1-75f6-4f6f-8994-36fe6f3b63f7" ;
		:name = "Attribute demonstration" ;
		:title = "Attribute demonstration" ;
data:

 x = -4, -2, 0, 2, 4 ;

 y = 50, 52, 54, 56, 58 ;

 alt = 50 ;

 time_instant = 27133200 ;

 time_instant_bounds =
  27133200, 27133200 ;

 time_counter = 27133200 ;

 time_counter_bounds =
  27133200, 27133200 ;

 forecast_reference_time = 27133200 ; 

 original_data =
  0, 2, 4, 6, 8,
  2, 4, 6, 8, 10,
  4, 6, 8, 10, 12,
  6, 8, 10, 12, 14,
  8, 10, 12, 14, 16 ;
}
